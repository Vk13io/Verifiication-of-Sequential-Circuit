
`include "uvm_macros.svh"
package tb_pkg;
 import uvm_pkg::*;
 `include "ring_sequence_item.sv"  
 `include "ring_sequence.sv"             
 `include "ring_sequencer.sv"           
 `include "ring_driver.sv"              
 `include "ring_monitor.sv"            
 `include "ring_agent.sv"                         
 `include "ring_scoreboard.sv"        
 `include "ring_env.sv"                
 `include "ring_test.sv"                

endpackage


